`timescale 1ns / 1ps

module Permuted_Choice2(LEFT_CIRCULAR_SHIFT1, RIGHT_CIRCULAR_SHIFT1, SUBKEY);

input [28 : 1] LEFT_CIRCULAR_SHIFT1;

input [28 : 1] RIGHT_CIRCULAR_SHIFT1;
output [48 : 1] SUBKEY;

wire [28 : 1] LEFT_CIRCULAR_SHIFT1;

wire [28 : 1] RIGHT_CIRCULAR_SHIFT1;
reg [48 : 1] SUBKEY;

wire [56 : 1] PERMUTATION2_INPUT;
 assign PERMUTATION2_INPUT = {LEFT_CIRCULAR_SHIFT1 , RIGHT_CIRCULAR_SHIFT1};
 always @ (PERMUTATION2_INPUT)
 begin
 SUBKEY[1] <= PERMUTATION2_INPUT[14];
 SUBKEY[2] <= PERMUTATION2_INPUT[17];
 SUBKEY[3] <= PERMUTATION2_INPUT[11];
 SUBKEY[4] <= PERMUTATION2_INPUT[24];
 SUBKEY[5] <= PERMUTATION2_INPUT[1];
 SUBKEY[6] <= PERMUTATION2_INPUT[5];
 SUBKEY[7] <= PERMUTATION2_INPUT[3];
 SUBKEY[8] <= PERMUTATION2_INPUT[28];
 SUBKEY[9] <= PERMUTATION2_INPUT[15];
 SUBKEY[10] <= PERMUTATION2_INPUT[6];
 SUBKEY[11] <= PERMUTATION2_INPUT[21];
 SUBKEY[12] <= PERMUTATION2_INPUT[10];
 SUBKEY[13] <= PERMUTATION2_INPUT[23];
 SUBKEY[14] <= PERMUTATION2_INPUT[19];
 SUBKEY[15] <= PERMUTATION2_INPUT[12];
 SUBKEY[16] <= PERMUTATION2_INPUT[4];
 SUBKEY[17] <= PERMUTATION2_INPUT[26];
 SUBKEY[18] <= PERMUTATION2_INPUT[8];
 SUBKEY[19] <= PERMUTATION2_INPUT[16];
 SUBKEY[20] <= PERMUTATION2_INPUT[7];
 SUBKEY[21] <= PERMUTATION2_INPUT[27];
 SUBKEY[22] <= PERMUTATION2_INPUT[20];
 SUBKEY[23] <= PERMUTATION2_INPUT[13];
 SUBKEY[24] <= PERMUTATION2_INPUT[2];
 SUBKEY[25] <= PERMUTATION2_INPUT[41];
 SUBKEY[26] <= PERMUTATION2_INPUT[52];
 SUBKEY[27] <= PERMUTATION2_INPUT[31];
 SUBKEY[28] <= PERMUTATION2_INPUT[37];
 SUBKEY[29] <= PERMUTATION2_INPUT[47];
 SUBKEY[30] <= PERMUTATION2_INPUT[55];
 SUBKEY[31] <= PERMUTATION2_INPUT[30];
 SUBKEY[32] <= PERMUTATION2_INPUT[40];
 SUBKEY[33] <= PERMUTATION2_INPUT[51];
 SUBKEY[34] <= PERMUTATION2_INPUT[45];
 SUBKEY[35] <= PERMUTATION2_INPUT[33];
 SUBKEY[36] <= PERMUTATION2_INPUT[48];
 SUBKEY[37] <= PERMUTATION2_INPUT[44];
 SUBKEY[38] <= PERMUTATION2_INPUT[49];
 SUBKEY[39] <= PERMUTATION2_INPUT[39];
SUBKEY[40] <= PERMUTATION2_INPUT[56];
SUBKEY[41] <= PERMUTATION2_INPUT[34];
SUBKEY[42] <= PERMUTATION2_INPUT[53];
SUBKEY[43] <= PERMUTATION2_INPUT[46];
SUBKEY[44] <= PERMUTATION2_INPUT[42];
SUBKEY[45] <= PERMUTATION2_INPUT[50];
SUBKEY[46] <= PERMUTATION2_INPUT[36];
SUBKEY[47] <= PERMUTATION2_INPUT[29];
SUBKEY[48] <= PERMUTATION2_INPUT[32];
end
endmodule
