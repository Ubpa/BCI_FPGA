`timescale 1ns / 1ps

module ip(PLAIN_TEXT, CHIP_SELECT_BAR, LEFT, RIGHT);
input CHIP_SELECT_BAR; 
input [64 : 1] PLAIN_TEXT ; 
output [32 : 1] LEFT;
output [32 : 1] RIGHT;
wire CHIP_SELECT_BAR;
wire [64 : 1] PLAIN_TEXT;
wire [32 : 1] LEFT;
wire [32 : 1] RIGHT;
 
reg [64 : 1] INITIAL_PERMUTATION_OUTPUT;
assign LEFT = INITIAL_PERMUTATION_OUTPUT[64 : 33];
assign RIGHT = INITIAL_PERMUTATION_OUTPUT[32 : 1];
always @ (*) 
begin
if(CHIP_SELECT_BAR == 0)
begin
INITIAL_PERMUTATION_OUTPUT [1] <= PLAIN_TEXT [58];
INITIAL_PERMUTATION_OUTPUT [2] <= PLAIN_TEXT [50];
INITIAL_PERMUTATION_OUTPUT [3] <= PLAIN_TEXT [42];
INITIAL_PERMUTATION_OUTPUT [4] <= PLAIN_TEXT [34];
INITIAL_PERMUTATION_OUTPUT [5] <= PLAIN_TEXT [26];
INITIAL_PERMUTATION_OUTPUT [6] <= PLAIN_TEXT [18];
INITIAL_PERMUTATION_OUTPUT [7] <= PLAIN_TEXT [10];
INITIAL_PERMUTATION_OUTPUT [8] <= PLAIN_TEXT [2];
INITIAL_PERMUTATION_OUTPUT [9] <= PLAIN_TEXT [60];
INITIAL_PERMUTATION_OUTPUT [10] <= PLAIN_TEXT [52];
INITIAL_PERMUTATION_OUTPUT [11] <= PLAIN_TEXT [44];
INITIAL_PERMUTATION_OUTPUT [12] <= PLAIN_TEXT [36];
INITIAL_PERMUTATION_OUTPUT [13] <= PLAIN_TEXT [28];
INITIAL_PERMUTATION_OUTPUT [14] <= PLAIN_TEXT [20];
INITIAL_PERMUTATION_OUTPUT [15] <= PLAIN_TEXT [12];
INITIAL_PERMUTATION_OUTPUT [16] <= PLAIN_TEXT [4];
INITIAL_PERMUTATION_OUTPUT [17] <= PLAIN_TEXT [62];
INITIAL_PERMUTATION_OUTPUT [18] <= PLAIN_TEXT [54];
INITIAL_PERMUTATION_OUTPUT [19] <= PLAIN_TEXT [46];
INITIAL_PERMUTATION_OUTPUT [20] <= PLAIN_TEXT [38];
INITIAL_PERMUTATION_OUTPUT [21] <= PLAIN_TEXT [30];
INITIAL_PERMUTATION_OUTPUT [22] <= PLAIN_TEXT [22];
INITIAL_PERMUTATION_OUTPUT [23] <= PLAIN_TEXT [14];
INITIAL_PERMUTATION_OUTPUT [24] <= PLAIN_TEXT [6];
INITIAL_PERMUTATION_OUTPUT [25] <= PLAIN_TEXT [64];
INITIAL_PERMUTATION_OUTPUT [26] <= PLAIN_TEXT [56];
INITIAL_PERMUTATION_OUTPUT [27] <= PLAIN_TEXT [48];
INITIAL_PERMUTATION_OUTPUT [28] <= PLAIN_TEXT [40];
INITIAL_PERMUTATION_OUTPUT [29] <= PLAIN_TEXT [32];
INITIAL_PERMUTATION_OUTPUT [30] <= PLAIN_TEXT [24];
INITIAL_PERMUTATION_OUTPUT [31] <= PLAIN_TEXT [16];
INITIAL_PERMUTATION_OUTPUT [32] <= PLAIN_TEXT [8];
INITIAL_PERMUTATION_OUTPUT [33] <= PLAIN_TEXT [57];
INITIAL_PERMUTATION_OUTPUT [34] <= PLAIN_TEXT [49];
INITIAL_PERMUTATION_OUTPUT [35] <= PLAIN_TEXT [41];
INITIAL_PERMUTATION_OUTPUT [36] <= PLAIN_TEXT [33];
INITIAL_PERMUTATION_OUTPUT [37] <= PLAIN_TEXT [25];
INITIAL_PERMUTATION_OUTPUT [38] <= PLAIN_TEXT [17];
INITIAL_PERMUTATION_OUTPUT [39] <= PLAIN_TEXT [9];
INITIAL_PERMUTATION_OUTPUT [40] <= PLAIN_TEXT [1];
INITIAL_PERMUTATION_OUTPUT [41] <= PLAIN_TEXT [59];
INITIAL_PERMUTATION_OUTPUT [42] <= PLAIN_TEXT [51];
INITIAL_PERMUTATION_OUTPUT [43] <= PLAIN_TEXT [43];
INITIAL_PERMUTATION_OUTPUT [44] <= PLAIN_TEXT [35];
INITIAL_PERMUTATION_OUTPUT [45] <= PLAIN_TEXT [27];
INITIAL_PERMUTATION_OUTPUT [46] <= PLAIN_TEXT [19];
INITIAL_PERMUTATION_OUTPUT [47] <= PLAIN_TEXT [11];
INITIAL_PERMUTATION_OUTPUT [48] <= PLAIN_TEXT [3];
INITIAL_PERMUTATION_OUTPUT [49] <= PLAIN_TEXT [61];
INITIAL_PERMUTATION_OUTPUT [50] <= PLAIN_TEXT [53];
INITIAL_PERMUTATION_OUTPUT [51] <= PLAIN_TEXT [45];
INITIAL_PERMUTATION_OUTPUT [52] <= PLAIN_TEXT [37];
INITIAL_PERMUTATION_OUTPUT [53] <= PLAIN_TEXT [29];
INITIAL_PERMUTATION_OUTPUT [54] <= PLAIN_TEXT [21];
INITIAL_PERMUTATION_OUTPUT [55] <= PLAIN_TEXT [13];
INITIAL_PERMUTATION_OUTPUT [56] <= PLAIN_TEXT [5];
INITIAL_PERMUTATION_OUTPUT [57] <= PLAIN_TEXT [63];
INITIAL_PERMUTATION_OUTPUT [58] <= PLAIN_TEXT [55];
INITIAL_PERMUTATION_OUTPUT [59] <= PLAIN_TEXT [47];
INITIAL_PERMUTATION_OUTPUT [60] <= PLAIN_TEXT [39];
INITIAL_PERMUTATION_OUTPUT [61] <= PLAIN_TEXT [31];
INITIAL_PERMUTATION_OUTPUT [62] <= PLAIN_TEXT [23];
INITIAL_PERMUTATION_OUTPUT [63] <= PLAIN_TEXT [15];
INITIAL_PERMUTATION_OUTPUT [64] <= PLAIN_TEXT [7];
end
else
begin
INITIAL_PERMUTATION_OUTPUT [64 : 1] <= 64'b0;
end
end
endmodule

